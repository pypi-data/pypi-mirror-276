// GENERATE INPLACE BEGIN fileheader() =========================================
//
// Module:     glbl.clk_gate
// Data Model: glbl.clk_gate.ClkGateMod
//
// GENERATE INPLACE END fileheader =============================================

// GENERATE INPLACE BEGIN header() =============================================
// GENERATE INPLACE END header =================================================

// GENERATE INPLACE BEGIN beginmod() ===========================================
module clk_gate ( // glbl.clk_gate.ClkGateMod
  input  wire  clk_i,
  output logic clk_o,
  input  wire  ena_i
);
// GENERATE INPLACE END beginmod ===============================================

    // GENERATE INPLACE BEGIN logic() ==========================================
    // GENERATE INPLACE END logic ==============================================

// GENERATE INPLACE BEGIN endmod() =============================================
endmodule // clk_gate
// GENERATE INPLACE END endmod =================================================

// GENERATE INPLACE BEGIN footer() =============================================
// GENERATE INPLACE END footer =================================================
